* RCA3040 CKT - RCA 3040 WIDEBAND AMPLIFIER.

.MODEL QNL NPN BF=80 RB=100 CJS=2p TF=0.3NS TR=6NS CJE=3PF CJC=2PF VAF=50

VIN 1 0 SIN (0 0.1 50MEG 0.5NS 0.0)
VCC 2 0 15.0
VEE 3 0 -15.0
RS1 30 1 1K
RS2 31 0 1K
R1 5 3 4.8K
R2 6 3 4.8K
R3 9 3 811
R4 8 3 2.17K
R5 8 0 820
R6 2 14 1.32K
R7 2 12 4.5K
R8 2 15 1.32K
R9 16 0 5.25K
R10 17 0 5.25K
Q1 2 30 5  QNL
Q2 2 31 6  QNL
Q3 10 5 7  QNL
Q4 11 6 7  QNL
Q5 14 12 10  QNL
Q6 15 12 11  QNL
Q7 12 12 13  QNL
Q8 13 13 0  QNL
Q9 7 8 9  QNL
Q10 2 15 16  QNL
Q11 2 14 17  QNL

*
*.PRINT TRAN V(1) V(16) V(17)
*.TRAN 0.5NS 200NS
*.OPTIONS LIMPTS=501
.END
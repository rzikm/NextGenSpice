SBDGATE CKT - SCHOTTKY-BARRIER TTL INVERTER

.MODEL D2 D(RS=15 CJO=0.2PF IS=5e-10 )
.MODEL QND NPN(BF=50 RB=70 RC=40 CJS=2PF TF=0.1NS TR=10NS
+ CJE=0.9PF CJC=1.5PF VJC=0.85 VAF=50)

VCC 23 0 5.0
VLOAD 26 0 5.0
VIN 1 0 PULSE 0.2 3.6 2NS 2NS 2NS 50NS

RS 1 2 50
RB1 23 3 15K
RB2 26 17 15K
RC1 4 5 60
RC2 6 9 30
RC3 16 15 10
RC4 18 19 60
RE1 7 8 600
RE2 20 21 600
RL1 23 10 8.75K
RL2 26 25 8K
RK 23 12 1K
RS2 24 15 50
Q1 4 3 2 QND
Q2 6 5 7 QND
Q3 16 7 0 QND
Q4 18 17 24 QND
Q5 22 19 20 QND
Q6 20 20 0 QND
QL2 25 25 22 QND
QE 12 10 13 QND
DC1 3 4 D2
DC2 5 6 D2
DC3 7 16 D2
DC4 17 18 D2
DC5 19 22 D2
DE1 8 0 D2
DE2 21 0 D2
D1 13 14 D2
D12 14 28 D2
D2 28 15 D2
DL 10 9 D2


*.TRAN 1NS 200NS
*.PRINT TRAN V(1) V(15) I(VCC)
.END

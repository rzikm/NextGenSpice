DIFPAIR CKT - SIMPLE DIFFERENTIAL PAIR
*
.MODEL QNL NPN(BF=80 RB=100 CJS=2PF TF=0.3NS TR=6NS CJE=3PF CJC=2PF VAF=50)
VIN 1 0 SIN(0.0 0.1 5MEG 5NS)
VCC 8 0 12
VEE 9 0 -12
Q1 4 2 6 QNL
Q2 5 3 6 QNL
RS1 1 2 1K
RS2 3 0 1K
RC1 4 8 10K
RC2 5 8 10K
Q3 6 7 9 QNL
Q4 7 7 9 QNL
RBIAS 7 8 20K

*.TRAN 5ns 500ns
*.PRINT TRAN V(1) V(4) V(5) 
.END

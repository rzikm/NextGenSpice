* ECL CKT - EMITTER COUPLED LOGIC INVERTER

VIN 1 0 PULSE(-1.0 -1.8 1NS 1NS 8NS 20NS)
VEE 8 0 -5.0
VREF 6 0 -1.4
Q1 3 2 4 QSTD
Q2 5 6 4 QSTD
Q3 0 5 7 QSTD
Q4 0 5 7 QSTD
RIN 1 2 50
RC1 0 3 120
RC2 0 5 135
RE 4 8 340
RTH1 7 8 125
RTH2 7 0 85
CLOAD 7 0 5P

.MODEL QSTD NPN IS=1E-16 BF=50 BR=0.1 RB=50 RC=10 TF=0.12N
+  TR=5N CJE=0.4P VJE=0.8 MJE=0.4 CJC=0.5P VJC=0.8 MJC=0.333
+  CJS=1P VAF=50

*.OPTIONS ABSTOL=1E-12 RELTOL=1E-5
*.TRAN 0.2NS 10NS
*.PRINT TRAN V(1) V(3) V(5) V(7) I(VIN)
.END

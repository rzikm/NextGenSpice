UA709 CKT - UA 709 OPERATIONAL AMPLIFIER
*
VIN 1 0 SIN 0 0.1 10K 2.5US 0
VCC 19 0 DC 15.0
VEE 20 0 DC -15.0
RS1 30 1 1K
RS2 31 0 1K
RF 30 18 100K
RCOMP 7 23 1.5K
CICOMP 23 2 5000PF
COCOMP 18 15 200PF

Q1 2 30 3  QNL
Q2 4 31 3  QNL
Q3 19 6 5  QNL
Q4 6 4 11  QNL
Q5 6 11 12  QNL
Q6 7 13 12  QNL
Q7 7 2 13  QNL
Q8 19 7 21  QNL
Q9 19 17 18  QNL
Q10 17 15 16  QNL
Q11 3 8 22  QNL
Q12 8 8 20  QNL
Q13 14 14 12  QNL
Q14 15 12 10  QPL
Q15 20 17 18  QPL
R1 5 2 25K
R2 5 4 25K
R3 22 20 2.4K
R4 8 9 18K
R5 9 12 3.6K
R6 11 14 3K
R7 19 6 10K
R8 19 7 10K
R9 9 10 10K
R10 10 18 30K
R11 19 17 20K
R12 15 16 10K
R13 16 20 75
R14 13 14 3K
R15 21 10 1K
.MODEL QNL NPN BF=80 RB=100 CJS=2p TF=0.3NS TR=6NS CJE=3PF CJC=2PF VAF=50
.MODEL QPL PNP BF=10 RB=20  TF=1NS   TR=20NS CJE=6PF CJC=4PF VAF=50
*
*.PRINT TRAN V(1) V(30) V(7) V(18)
*.TRAN 2.0US 250US
*.OPTIONS RELTOL=1E-5
.END
